module int2fp (
    input  [31:0] A,
    output reg [31:0] B
);

    reg [31:0] abs;
    reg        sign;
    reg [22:0] mout;      // mantissa
    reg [7:0]  eout;      // exponent
    reg [7:0]  num_zeros;

    always @(*) begin
        // Calcula o valor absoluto e sinal
        abs  = (A[31]) ? (~A + 32'd1) : A;

        if (abs[30:0] == 0) begin
            // Valor zero
            eout       = 8'd0;
            mout       = 23'd0;
            sign       = 1'b0;
            num_zeros  = 8'd0;
        end 
        else begin
            // Determina o número de zeros à esquerda (normalização)
            casez (abs[30:0])
                31'b1???????????????????????????????: num_zeros = 8'd0;
                31'b01??????????????????????????????: num_zeros = 8'd1;
                31'b001?????????????????????????????: num_zeros = 8'd2;
                31'b0001????????????????????????????: num_zeros = 8'd3;
                31'b00001???????????????????????????: num_zeros = 8'd4;
                31'b000001??????????????????????????: num_zeros = 8'd5;
                31'b0000001?????????????????????????: num_zeros = 8'd6;
                31'b00000001????????????????????????: num_zeros = 8'd7;
                31'b000000001???????????????????????: num_zeros = 8'd8;
                31'b0000000001??????????????????????: num_zeros = 8'd9;
                31'b00000000001?????????????????????: num_zeros = 8'd10;
                31'b000000000001????????????????????: num_zeros = 8'd11;
                31'b0000000000001???????????????????: num_zeros = 8'd12;
                31'b00000000000001??????????????????: num_zeros = 8'd13;
                31'b000000000000001?????????????????: num_zeros = 8'd14;
                31'b0000000000000001????????????????: num_zeros = 8'd15;
                31'b00000000000000001???????????????: num_zeros = 8'd16;
                31'b000000000000000001??????????????: num_zeros = 8'd17;
                31'b0000000000000000001?????????????: num_zeros = 8'd18;
                31'b00000000000000000001????????????: num_zeros = 8'd19;
                31'b000000000000000000001???????????: num_zeros = 8'd20;
                31'b0000000000000000000001??????????: num_zeros = 8'd21;
                31'b00000000000000000000001?????????: num_zeros = 8'd22;
                31'b000000000000000000000001????????: num_zeros = 8'd23;
                31'b0000000000000000000000001???????: num_zeros = 8'd24;
                31'b00000000000000000000000001??????: num_zeros = 8'd25;
                31'b000000000000000000000000001?????: num_zeros = 8'd26;
                31'b0000000000000000000000000001????: num_zeros = 8'd27;
                31'b00000000000000000000000000001???: num_zeros = 8'd28;
                31'b000000000000000000000000000001??: num_zeros = 8'd29;
                31'b0000000000000000000000000000001?: num_zeros = 8'd30;
                31'b00000000000000000000000000000001: num_zeros = 8'd31;
                default: num_zeros = 8'd31;
            endcase

            // Normaliza e calcula expoente
            mout = (abs[30:0] << num_zeros) >> 7;
            eout = 8'd157 - num_zeros;  // 127 + 30 = 157
            sign = A[31];
        end

        // Monta o número em ponto flutuante IEEE 754
        B = {sign, eout, mout};
    end

endmodule
